../../../../modelsimPatch/vhdl/simulationPkg/simulationPkg.vhd