library ieee;
use ieee.std_logic_1164.all;

entity switchTb is
	-- Testbench has no input and output signals!
end switchTb;

architecture testbench of switchTb is
begin
	
	
	
end architecture testbench;
